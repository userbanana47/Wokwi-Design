// Copyright 2025 Michael Schurz
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE−2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

//`timescale 1ns / 1ps

module button_pulse(
	input wire clk,
	input wire reset,
	input wire btn,
	output reg pulse
);
	reg last_btn;
	always @(posedge clk or posedge reset) begin
		if (reset) begin
			pulse <= 0;
			last_btn <= 0;
		end else begin
			last_btn <= btn;
			pulse <= btn && ~last_btn;
		end
	end
endmodule
